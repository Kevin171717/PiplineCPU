module shifter(input [31:0] dataIn, input [4:0] amount, input select, output [31:0] dataOut);
    wire[4:0] shift;
    assign shift = select ? amount : 5'b00000;
    wire [31:0] stage0, stage1, stage2, stage3, stage4;

    assign stage0[0]  = shift[0] ? 1'b0       : dataIn[0];
    assign stage0[1]  = shift[0] ? dataIn[0]  : dataIn[1];
    assign stage0[2]  = shift[0] ? dataIn[1]  : dataIn[2];
    assign stage0[3]  = shift[0] ? dataIn[2]  : dataIn[3];
    assign stage0[4]  = shift[0] ? dataIn[3]  : dataIn[4];
    assign stage0[5]  = shift[0] ? dataIn[4]  : dataIn[5];
    assign stage0[6]  = shift[0] ? dataIn[5]  : dataIn[6];
    assign stage0[7]  = shift[0] ? dataIn[6]  : dataIn[7];
    assign stage0[8]  = shift[0] ? dataIn[7]  : dataIn[8];
    assign stage0[9]  = shift[0] ? dataIn[8]  : dataIn[9];
    assign stage0[10] = shift[0] ? dataIn[9]  : dataIn[10];
    assign stage0[11] = shift[0] ? dataIn[10] : dataIn[11];
    assign stage0[12] = shift[0] ? dataIn[11] : dataIn[12];
    assign stage0[13] = shift[0] ? dataIn[12] : dataIn[13];
    assign stage0[14] = shift[0] ? dataIn[13] : dataIn[14];
    assign stage0[15] = shift[0] ? dataIn[14] : dataIn[15];
    assign stage0[16] = shift[0] ? dataIn[15] : dataIn[16];
    assign stage0[17] = shift[0] ? dataIn[16] : dataIn[17];
    assign stage0[18] = shift[0] ? dataIn[17] : dataIn[18];
    assign stage0[19] = shift[0] ? dataIn[18] : dataIn[19];
    assign stage0[20] = shift[0] ? dataIn[19] : dataIn[20];
    assign stage0[21] = shift[0] ? dataIn[20] : dataIn[21];
    assign stage0[22] = shift[0] ? dataIn[21] : dataIn[22];
    assign stage0[23] = shift[0] ? dataIn[22] : dataIn[23];
    assign stage0[24] = shift[0] ? dataIn[23] : dataIn[24];
    assign stage0[25] = shift[0] ? dataIn[24] : dataIn[25];
    assign stage0[26] = shift[0] ? dataIn[25] : dataIn[26];
    assign stage0[27] = shift[0] ? dataIn[26] : dataIn[27];
    assign stage0[28] = shift[0] ? dataIn[27] : dataIn[28];
    assign stage0[29] = shift[0] ? dataIn[28] : dataIn[29];
    assign stage0[30] = shift[0] ? dataIn[29] : dataIn[30];
    assign stage0[31] = shift[0] ? dataIn[30] : dataIn[31];


    assign stage1[0]  = shift[1] ? 1'b0       : stage0[0];
    assign stage1[1]  = shift[1] ? 1'b0       : stage0[1];
    assign stage1[2]  = shift[1] ? stage0[0]  : stage0[2];
    assign stage1[3]  = shift[1] ? stage0[1]  : stage0[3];
    assign stage1[4]  = shift[1] ? stage0[2]  : stage0[4];
    assign stage1[5]  = shift[1] ? stage0[3]  : stage0[5];
    assign stage1[6]  = shift[1] ? stage0[4]  : stage0[6];
    assign stage1[7]  = shift[1] ? stage0[5]  : stage0[7];
    assign stage1[8]  = shift[1] ? stage0[6]  : stage0[8];
    assign stage1[9]  = shift[1] ? stage0[7]  : stage0[9];
    assign stage1[10] = shift[1] ? stage0[8]  : stage0[10];
    assign stage1[11] = shift[1] ? stage0[9]  : stage0[11];
    assign stage1[12] = shift[1] ? stage0[10] : stage0[12];
    assign stage1[13] = shift[1] ? stage0[11] : stage0[13];
    assign stage1[14] = shift[1] ? stage0[12] : stage0[14];
    assign stage1[15] = shift[1] ? stage0[13] : stage0[15];
    assign stage1[16] = shift[1] ? stage0[14] : stage0[16];
    assign stage1[17] = shift[1] ? stage0[15] : stage0[17];
    assign stage1[18] = shift[1] ? stage0[16] : stage0[18];
    assign stage1[19] = shift[1] ? stage0[17] : stage0[19];
    assign stage1[20] = shift[1] ? stage0[18] : stage0[20];
    assign stage1[21] = shift[1] ? stage0[19] : stage0[21];
    assign stage1[22] = shift[1] ? stage0[20] : stage0[22];
    assign stage1[23] = shift[1] ? stage0[21] : stage0[23];
    assign stage1[24] = shift[1] ? stage0[22] : stage0[24];
    assign stage1[25] = shift[1] ? stage0[23] : stage0[25];
    assign stage1[26] = shift[1] ? stage0[24] : stage0[26];
    assign stage1[27] = shift[1] ? stage0[25] : stage0[27];
    assign stage1[28] = shift[1] ? stage0[26] : stage0[28];
    assign stage1[29] = shift[1] ? stage0[27] : stage0[29];
    assign stage1[30] = shift[1] ? stage0[28] : stage0[30];
    assign stage1[31] = shift[1] ? stage0[29] : stage0[31];


    assign stage2[0]  = shift[2] ? 1'b0 : stage1[0];
    assign stage2[1]  = shift[2] ? 1'b0 : stage1[1];
    assign stage2[2]  = shift[2] ? 1'b0 : stage1[2];
    assign stage2[3]  = shift[2] ? 1'b0 : stage1[3];
    assign stage2[4]  = shift[2] ? stage1[0] : stage1[4];
    assign stage2[5]  = shift[2] ? stage1[1] : stage1[5];
    assign stage2[6]  = shift[2] ? stage1[2] : stage1[6];
    assign stage2[7]  = shift[2] ? stage1[3] : stage1[7];
    assign stage2[8]  = shift[2] ? stage1[4] : stage1[8];
    assign stage2[9]  = shift[2] ? stage1[5] : stage1[9];
    assign stage2[10] = shift[2] ? stage1[6] : stage1[10];
    assign stage2[11] = shift[2] ? stage1[7] : stage1[11];
    assign stage2[12] = shift[2] ? stage1[8] : stage1[12];
    assign stage2[13] = shift[2] ? stage1[9] : stage1[13];
    assign stage2[14] = shift[2] ? stage1[10] : stage1[14];
    assign stage2[15] = shift[2] ? stage1[11] : stage1[15];
    assign stage2[16] = shift[2] ? stage1[12] : stage1[16];
    assign stage2[17] = shift[2] ? stage1[13] : stage1[17];
    assign stage2[18] = shift[2] ? stage1[14] : stage1[18];
    assign stage2[19] = shift[2] ? stage1[15] : stage1[19];
    assign stage2[20] = shift[2] ? stage1[16] : stage1[20];
    assign stage2[21] = shift[2] ? stage1[17] : stage1[21];
    assign stage2[22] = shift[2] ? stage1[18] : stage1[22];
    assign stage2[23] = shift[2] ? stage1[19] : stage1[23];
    assign stage2[24] = shift[2] ? stage1[20] : stage1[24];
    assign stage2[25] = shift[2] ? stage1[21] : stage1[25];
    assign stage2[26] = shift[2] ? stage1[22] : stage1[26];
    assign stage2[27] = shift[2] ? stage1[23] : stage1[27];
    assign stage2[28] = shift[2] ? stage1[24] : stage1[28];
    assign stage2[29] = shift[2] ? stage1[25] : stage1[29];
    assign stage2[30] = shift[2] ? stage1[26] : stage1[30];
    assign stage2[31] = shift[2] ? stage1[27] : stage1[31];


    assign stage3[0]  = shift[3] ? 1'b0 : stage2[0];
    assign stage3[1]  = shift[3] ? 1'b0 : stage2[1];
    assign stage3[2]  = shift[3] ? 1'b0 : stage2[2];
    assign stage3[3]  = shift[3] ? 1'b0 : stage2[3];
    assign stage3[4]  = shift[3] ? 1'b0 : stage2[4];
    assign stage3[5]  = shift[3] ? 1'b0 : stage2[5];
    assign stage3[6]  = shift[3] ? 1'b0 : stage2[6];
    assign stage3[7]  = shift[3] ? 1'b0 : stage2[7];
    assign stage3[8]  = shift[3] ? stage2[0] : stage2[8];
    assign stage3[9]  = shift[3] ? stage2[1] : stage2[9];
    assign stage3[10] = shift[3] ? stage2[2] : stage2[10];
    assign stage3[11] = shift[3] ? stage2[3] : stage2[11];
    assign stage3[12] = shift[3] ? stage2[4] : stage2[12];
    assign stage3[13] = shift[3] ? stage2[5] : stage2[13];
    assign stage3[14] = shift[3] ? stage2[6] : stage2[14];
    assign stage3[15] = shift[3] ? stage2[7] : stage2[15];
    assign stage3[16] = shift[3] ? stage2[8] : stage2[16];
    assign stage3[17] = shift[3] ? stage2[9] : stage2[17];
    assign stage3[18] = shift[3] ? stage2[10] : stage2[18];
    assign stage3[19] = shift[3] ? stage2[11] : stage2[19];
    assign stage3[20] = shift[3] ? stage2[12] : stage2[20];
    assign stage3[21] = shift[3] ? stage2[13] : stage2[21];
    assign stage3[22] = shift[3] ? stage2[14] : stage2[22];
    assign stage3[23] = shift[3] ? stage2[15] : stage2[23];
    assign stage3[24] = shift[3] ? stage2[16] : stage2[24];
    assign stage3[25] = shift[3] ? stage2[17] : stage2[25];
    assign stage3[26] = shift[3] ? stage2[18] : stage2[26];
    assign stage3[27] = shift[3] ? stage2[19] : stage2[27];
    assign stage3[28] = shift[3] ? stage2[20] : stage2[28];
    assign stage3[29] = shift[3] ? stage2[21] : stage2[29];
    assign stage3[30] = shift[3] ? stage2[22] : stage2[30];
    assign stage3[31] = shift[3] ? stage2[23] : stage2[31];


    assign stage4[0]  = shift[4] ? 1'b0 : stage3[0];
    assign stage4[1]  = shift[4] ? 1'b0 : stage3[1];
    assign stage4[2]  = shift[4] ? 1'b0 : stage3[2];
    assign stage4[3]  = shift[4] ? 1'b0 : stage3[3];
    assign stage4[4]  = shift[4] ? 1'b0 : stage3[4];
    assign stage4[5]  = shift[4] ? 1'b0 : stage3[5];
    assign stage4[6]  = shift[4] ? 1'b0 : stage3[6];
    assign stage4[7]  = shift[4] ? 1'b0 : stage3[7];
    assign stage4[8]  = shift[4] ? 1'b0 : stage3[8];
    assign stage4[9]  = shift[4] ? 1'b0 : stage3[9];
    assign stage4[10] = shift[4] ? 1'b0 : stage3[10];
    assign stage4[11] = shift[4] ? 1'b0 : stage3[11];
    assign stage4[12] = shift[4] ? 1'b0 : stage3[12];
    assign stage4[13] = shift[4] ? 1'b0 : stage3[13];
    assign stage4[14] = shift[4] ? 1'b0 : stage3[14];
    assign stage4[15] = shift[4] ? 1'b0 : stage3[15];
    assign stage4[16] = shift[4] ? stage3[0] : stage3[16];
    assign stage4[17] = shift[4] ? stage3[1] : stage3[17];
    assign stage4[18] = shift[4] ? stage3[2] : stage3[18];
    assign stage4[19] = shift[4] ? stage3[3] : stage3[19];
    assign stage4[20] = shift[4] ? stage3[4] : stage3[20];
    assign stage4[21] = shift[4] ? stage3[5] : stage3[21];
    assign stage4[22] = shift[4] ? stage3[6] : stage3[22];
    assign stage4[23] = shift[4] ? stage3[7] : stage3[23];
    assign stage4[24] = shift[4] ? stage3[8] : stage3[24];
    assign stage4[25] = shift[4] ? stage3[9] : stage3[25];
    assign stage4[26] = shift[4] ? stage3[10] : stage3[26];
    assign stage4[27] = shift[4] ? stage3[11] : stage3[27];
    assign stage4[28] = shift[4] ? stage3[12] : stage3[28];
    assign stage4[29] = shift[4] ? stage3[13] : stage3[29];
    assign stage4[30] = shift[4] ? stage3[14] : stage3[30];
    assign stage4[31] = shift[4] ? stage3[15] : stage3[31];


    assign dataOut = stage4;
endmodule