module branchMUX();
endmodule